`timescale 1ns / 1ps;

module TestALU();
    reg [5:0] a;
    reg [5:0] b;
    reg [2:0] op;
    wire [5:0] res;
    wire err;
    
    ALU CUT (a, b, op, res, err);
    
    // Result range = [-32, 31]

    initial begin
        // Addition tests (opcode 0)
        op = 3'b000;
        a = 6'b001001; b = 6'b001010; #10;  // 9 + 10 = 19
        b = 6'b111100; #10;  // 9 + (-4) = 5
        b = 6'b110101; #10;  // 9 + (-11) = -2 
        a = 6'b010000; b = 6'b010111; #10;  // 16 + 23 = 39 (overflow)
        a = 6'b111000; b = 6'b111100; #10;  // (-8) + (-4) = -12
        // Subtraction tests (opcode 1)
        op = 3'b001;
        a = 6'b001010; b = 6'b001001; #10;  // 10 - 9 = 1
        a = 6'b001001; b = 6'b001010; #10;  // 9 - 10 = -1 - TODO: fix
        a = 6'b001001; b = 6'b111100; #10;  // 9 - (-4) = 13
        a = 6'b111100; b = 6'b001001; #10;  // (-4) - 9 = -13
        a = 6'b111100; b = 6'b110111; #10;  // (-4) - (-9) = 5
        a = 6'b110000; b = 6'b010111; #10;  // (-16) - 23 = -39 (underflow)
        // Decrement tests (opcode 2)
        op = 3'b010;
        a = 6'b001010; #10;  // 10 - 1 = 9
        a = 6'b111111; #10;  // 1 - 1 = 0
        a = 6'b000000; #10;  // 0 - 1 = -1
        a = 6'b110110; #10  // -10 - 1 = -11
        a = 6'b100000; #10  // -32 - 1 = -33 (overflow)
        // Increment tests (opcode 3)
        op = 3'b011;
        a = 6'b001010; #10;  // 10 + 1 = 11
        a = 6'b000000; #10;  // 0 + 1 = 1
        a = 6'b111111; #10;  // -1 + 1 = 0
        a = 6'b110110; #10;  // -10 + 1 = 9
        a = 6'b011111; #10;  // 31 + 1 = 32 (overflow)
        // Bitwise NOT tests (opcode 4)
        op = 3'b100;
        a = 6'b000000; #10;  // ~000000 = 111111
        a = 6'b111111; #10;  // ~111111 = 000000
        a = 6'b000111; #10;  // ~000111 = 111000
        // Bitwise AND tests (opcode 5)
        op = 3'b101;
        a = 6'b000000; b = 6'b111111; #10;  // 000000 & 111111 = 000000
        a = 6'b111111; b = 6'b000000; #10;  // 111111 & 000000 = 000000
        a = 6'b000111; b = 6'b111111; #10;  // 000111 & 111111 = 000111
        a = 6'b000111; b = 6'b000000; #10;  // 000111 & 000000 = 000000
        // Bitwise OR tests (opcode 6)
        op = 3'b110;
        a = 6'b000000; b = 6'b111111; #10;  // 000000 | 111111 = 111111
        a = 6'b111111; b = 6'b000000; #10;  // 111111 | 000000 = 111111
        a = 6'b000111; b = 6'b111111; #10;  // 000111 | 111111 = 111111
        a = 6'b000111; b = 6'b000000; #10;  // 000111 | 000000 = 000111
        // Bitwise XOR tests (opcode 7)
        op = 3'b111;
        a = 6'b000000; b = 6'b111111; #10;  // 000000 ^ 111111 = 111111
        a = 6'b111111; b = 6'b000000; #10;  // 111111 ^ 000000 = 111111
        a = 6'b000111; b = 6'b111111; #10;  // 000111 ^ 111111 = 000000
        a = 6'b000111; b = 6'b000000; #10;  // 000111 ^ 000000 = 000111
        $stop;
    end
endmodule
